module nimidecode(
input wire [31:0]ins,
input wire [1:0]msu,
input wire [5:0]statu_biu,
