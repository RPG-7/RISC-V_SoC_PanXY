module PERI_MUX
	(
		input HRESETn,
		input HCLK,
		input [31:0]PERISEL,
		output [31:0]PERIDATAR,
		output PERIREADY,
		input [31:0]PERIDATA0,
		input [31:0]PERIDATA1,
		input [31:0]PERIDATA2,
		input [31:0]PERIDATA3,
		input [31:0]PERIDATA4,
		input [31:0]PERIDATA5,
		input [31:0]PERIDATA6,
		input [31:0]PERIDATA7,
		
		input PERIREADY0,
		input PERIREADY1,
		input PERIREADY2,
		input PERIREADY3,
		input PERIREADY4,
		input PERIREADY5,
		input PERIREADY6,
		input PERIREADY7
	);
	reg[4:0]SLAVESEL;
	wire[4:0]SRDCO;
	always @(posedge HCLK or negedge HRESETn)
	begin
		if(!HRESETn)
			SLAVESEL<=1'b0;
		else
			SLAVESEL<=(PERIREADY)?(SRDCO):SLAVESEL;
	end
	assign SRDCO=(
		{5{PERISEL==	32'b10000000000000000000000000000000	}}&31|
		{5{PERISEL==	32'b01000000000000000000000000000000	}}&30|
		{5{PERISEL==	32'b00100000000000000000000000000000	}}&29|
		{5{PERISEL==	32'b00010000000000000000000000000000	}}&28|
		{5{PERISEL==	32'b00001000000000000000000000000000	}}&27|
		{5{PERISEL==	32'b00000100000000000000000000000000	}}&26|
		{5{PERISEL==	32'b00000010000000000000000000000000	}}&25|
		{5{PERISEL==	32'b00000001000000000000000000000000	}}&24|
		{5{PERISEL==	32'b00000000100000000000000000000000	}}&23|
		{5{PERISEL==	32'b00000000010000000000000000000000	}}&22|
		{5{PERISEL==	32'b00000000001000000000000000000000	}}&21|
		{5{PERISEL==	32'b00000000000100000000000000000000	}}&20|
		{5{PERISEL==	32'b00000000000010000000000000000000	}}&19|
		{5{PERISEL==	32'b00000000000001000000000000000000	}}&18|
		{5{PERISEL==	32'b00000000000000100000000000000000	}}&17|
		{5{PERISEL==	32'b00000000000000010000000000000000	}}&16|
		{5{PERISEL==	32'b00000000000000001000000000000000	}}&15|
		{5{PERISEL==	32'b00000000000000000100000000000000	}}&14|
		{5{PERISEL==	32'b00000000000000000010000000000000	}}&13|
		{5{PERISEL==	32'b00000000000000000001000000000000	}}&12|
		{5{PERISEL==	32'b00000000000000000000100000000000	}}&11|
		{5{PERISEL==	32'b00000000000000000000010000000000	}}&10|
		{5{PERISEL==	32'b00000000000000000000001000000000	}}&9|
		{5{PERISEL==	32'b00000000000000000000000100000000	}}&8|
		{5{PERISEL==	32'b00000000000000000000000010000000	}}&7|
		{5{PERISEL==	32'b00000000000000000000000001000000	}}&6|
		{5{PERISEL==	32'b00000000000000000000000000100000	}}&5|
		{5{PERISEL==	32'b00000000000000000000000000010000	}}&4|
		{5{PERISEL==	32'b00000000000000000000000000001000	}}&3|
		{5{PERISEL==	32'b00000000000000000000000000000100	}}&2|
		{5{PERISEL==	32'b00000000000000000000000000000010	}}&1|
		32'h0);
	
	assign PERIDATAR=(
	({32{SRDCO==1}}&PERIDATA0)|
	({32{SRDCO==2}}&PERIDATA1)|
	({32{SRDCO==3}}&PERIDATA2)|
	({32{SRDCO==4}}&PERIDATA3)|
	({32{SRDCO==5}}&PERIDATA4)|
	({32{SRDCO==6}}&PERIDATA5)|
	({32{SRDCO==7}}&PERIDATA6)|
	({32{SRDCO==8}}&PERIDATA7)|
	32'b0
	);
	
	assign PERIREADY=
	((SRDCO==0)|
	((SRDCO==1)&PERIREADY0)|
	((SRDCO==2)&PERIREADY1)|
	((SRDCO==3)&PERIREADY2)|
	((SRDCO==4)&PERIREADY3)|
	((SRDCO==5)&PERIREADY4)|
	((SRDCO==6)&PERIREADY5)|
	((SRDCO==7)&PERIREADY6)|
	((SRDCO==8)&PERIREADY7));
	
	
	
	
endmodule